module pipeline
(
    
)