module fetch_stage(
    input [31:0]PC_in,
    input [31:0]instruction_in,
    input instruction_valid,
    input clk,
    input resetn,
    output reg PC_out,
    output reg instruction_out,
    output instruction_received,
    output instruction_enable
);

endmodule;