module pipe_reg(
    input clk,
    input resetn
);
    reg [31:0] PC;
    reg [31:0] inst;
endmodule;